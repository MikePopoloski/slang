module m;
    libmod lm();
endmodule

module n(I.m im);
endmodule

`define SOME_DEF
