package type_forward_a_pkg;
  typedef type_base_pkg::foo_t foo_t;
endpackage
