"system stuff!"