.WIDTH(WIDTH),
