`define SOMETHING 1337