/* hello */
`include "local.svh"
`include "nested/file.svh"
`include "../data/nested/file.svh"