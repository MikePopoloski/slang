package dup_pkg;
endpackage

package dup_pkg;
endpackage

module top;
endmodule