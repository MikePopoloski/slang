module Foo();

endmodule

module Bar();

    Foo f();

endmodule
