.WIDTH (WIDTH),
.ENABLE(ENABLE)
