`define FOO(a) logic [2:0] b = a
