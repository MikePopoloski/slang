module n;
    m m1();
    int `ID(foo) = 1;
endmodule
