package consts_pkg;
  localparam int unsigned WIDTH = 48;
  localparam int unsigned DEPTH = 16;
endpackage
