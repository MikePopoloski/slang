`begin_keywords "1800-2012"

`include "another_systemverilog.sv"

`end_keywords

module t();

  wire do;

endmodule
