`pragma once
`include "local.svh"