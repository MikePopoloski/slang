package type_forward_b_pkg;
  typedef type_base_pkg::foo_t foo_t;
endpackage
