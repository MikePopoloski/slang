module m;
    int i = $foo;
endmodule
