`include "macro.svh"

module other;
    `FOO(1);
endmodule
