`define BAR `__FILE__
`define FOO `BAR
