`pragma protect data_block
abcd
