package pkg;
    localparam int bar = 42;

    class C; endclass
endpackage
