`include "another_systemverilog.sv"

module t();

  wire do;

endmodule
