`include "nested_local.svh"
`include "nonexistent.svh"
