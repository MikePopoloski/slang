package multihop_mid_pkg;
  import consts_pkg::*;
  // First hop forwards WIDTH to match consts_pkg exactly.
  localparam int unsigned WIDTH = consts_pkg::WIDTH;
endpackage
