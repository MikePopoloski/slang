module main;
    initial begin
    	$display("Something: %d", `SOMETHING);
    end
endmodule