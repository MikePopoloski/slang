package explicit_import_pkg;
  // Re-export WIDTH purely via an explicit import of the original symbol.
  import consts_pkg::WIDTH;
endpackage
