package type_base_pkg;
  typedef logic [7:0] foo_t;
endpackage
