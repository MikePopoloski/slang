module top;
    mod1 m();
endmodule
