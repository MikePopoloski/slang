parameter int WIDTH  = 8,
parameter bit ENABLE = 1
