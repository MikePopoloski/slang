.ENABLE(ENABLE),
