// Just a test string
"test string"
