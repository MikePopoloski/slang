module m1();

    wire a;

    always_comb begin
        $display(a);
    end

endmodule
