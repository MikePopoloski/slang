module simple;
endmodule
