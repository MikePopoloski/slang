module m;
    libmod lm();
endmodule
