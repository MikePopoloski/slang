module k;
    logic [3:0] a;
    logic [2:0] b = a;
endmodule
