module m;
    libmod lm();
endmodule

`define SOME_DEF
