`include "infinite_chain.svh"
