"test string"
