`include "nested/macro.svh"

module m;
    logic [3:0] a;
    `FOO(a);
endmodule
