`include "file_defn.svh"
`FOO
