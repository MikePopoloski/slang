parameter p = 1;
