"test string"