module module1
#(
    parameter int P1 = 4,
    parameter int P2 = 5
)
(
    input  logic [P1-1:0]   in1,
    input  logic [P2-1:0]   in2,
    input  logic [3:0]      in3,

    output logic [P1-1:0]   out1,
    output logic [P1-1:0]   out2,
    output logic [P1-1:0]   out3
);

    always_comb out1 = in1;

    always_comb begin
        out2 = in2;
        out3 = in3;
    end

    logic [7:0] arr1 [2 * $bits(out2)];

    typedef struct {
        logic [$bits(arr1[0]):0] f1;
        logic [$bits(arr1[1]):0] f2;
    } type1;

    type1 x;

endmodule
