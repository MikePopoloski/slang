"system stuff!"
